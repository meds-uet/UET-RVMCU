`ifndef VERILATOR
`include "../defines/gpio_defs.svh"
`else
`include "gpio_defs.svh"
`endif
